-------------------------------------------------------------------------------
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: XpmL1Router
-- 
-- Note: Common-to-XpmApp interface defined here (see URL below)
--       https://confluence.slac.stanford.edu/x/rLyMCw
-------------------------------------------------------------------------------
-- This file is part of 'L2SI Core'. It is subject to
-- the license terms in the LICENSE.txt file found in the top-level directory
-- of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'L2SI Core', including this file, may be
-- copied, modified, propagated, or distributed except according to the terms
-- contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiStreamPkg.all;

library l2si_core;
use l2si_core.XpmPkg.all;

entity XpmL1Router is
   generic (
      TPD_G       : time         := 1 ns;
      NUM_LINKS_G : integer      := 1 );
   port (
     clk            : in  sl;
     rst            : in  sl;
     l1FeedbacksIn  : in  XpmL1FeedbackArray(NUM_LINKS_G-1 downto 0);
     l1InAcks       : out slv               (NUM_LINKS_G-1 downto 0);
     l1FeedbacksOut : out XpmL1FeedbackArray(XPM_PARTITIONS_C downto 0);
     l1OutAcks      : in  slv               (XPM_PARTITIONS_C downto 0) );
end XpmL1Router;

architecture top_level_app of XpmL1Router is

begin
   l1InAcks       <= (others=>'1');
   l1FeedbacksOut <= (others=>XPM_L1_FEEDBACK_INIT_C);
end top_level_app;
