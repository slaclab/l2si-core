
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

package XpmOpts is

  constant TPGMINI_C : boolean := false;
  
end XpmOpts;
