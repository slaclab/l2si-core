
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use work.StdRtlPkg.all;

package FpgaTypePkg is

  constant CPSW_TARBALL_ADDR_C : slv(31 downto 0) := (others=>'0');
  
end FpgaTypePkg;
