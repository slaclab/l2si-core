weaver@pslab01.slac.stanford.edu.55856:1498499329