------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : XpmReg.vhd
-- Author     : Matt Weaver
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2015-12-14
-- Last update: 2017-03-31
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Software programmable register interface
-------------------------------------------------------------------------------
-- This file is part of 'LCLS2 XPM Core'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'LCLS2 XPM Core', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

use work.StdRtlPkg.all;
use work.AxiLitePkg.all;
use work.AxiStreamPkg.all;
use work.SsiPkg.all;
use work.AmcCarrierPkg.all;  -- ETH_AXIS_CONFIG_C
use work.XpmPkg.all;

entity XpmReg is
   port (
      axilClk          : in  sl;
      axilRst          : in  sl;
      axilUpdate       : out slv(NPartitions-1 downto 0);
      axilWriteMaster  : in  AxiLiteWriteMasterType;  
      axilWriteSlave   : out AxiLiteWriteSlaveType;  
      axilReadMaster   : in  AxiLiteReadMasterType;  
      axilReadSlave    : out AxiLiteReadSlaveType;
      -- Application Debug Interface (sysclk domain)
      ibDebugMaster    : in  AxiStreamMasterType;
      ibDebugSlave     : out AxiStreamSlaveType;
      --
      staClk           : in  sl;
      pllStatus        : in  XpmPllStatusArray(NAmcs-1 downto 0);
      status           : in  XpmStatusType;
      config           : out XpmConfigType;
      dbgChan          : out slv(4 downto 0) );
end XpmReg;

architecture rtl of XpmReg is

  type StateType is (IDLE_S, READING_S);
  
  type RegType is record
    state          : StateType;
    tagSlave       : AxiStreamSlaveType;
    load           : sl;
    config         : XpmConfigType;
    partition      : slv(3 downto 0);
    link           : slv(4 downto 0);
    amc            : slv(0 downto 0);
    inhibit        : slv(1 downto 0);
    linkCfg        : XpmLinkConfigType;
    linkStat       : XpmLinkStatusType;
    partitionCfg   : XpmPartitionConfigType;
    partitionStat  : XpmPartitionStatusType;
    pllCfg         : XpmPllConfigType;
    pllStat        : XpmPllStatusType;
    inhibitCfg     : XpmInhibitConfigType;
    axilReadSlave  : AxiLiteReadSlaveType;
    axilWriteSlave : AxiLiteWriteSlaveType;
    axilRdEn       : slv(NPartitions-1 downto 0);
    linkDebug      : slv(4 downto 0);
    tagStream      : sl;
    anaWrCount     : Slv32Array(NPartitions-1 downto 0);
  end record RegType;

  constant REG_INIT_C : RegType := (
    state          => IDLE_S,
    tagSlave       => AXI_STREAM_SLAVE_INIT_C,
    load           => '1',
    config         => XPM_CONFIG_INIT_C,
    partition      => (others=>'0'),
    link           => (others=>'0'),
    amc            => (others=>'0'),
    inhibit        => (others=>'0'),
    linkCfg        => XPM_LINK_CONFIG_INIT_C,
    linkStat       => XPM_LINK_STATUS_INIT_C,
    partitionCfg   => XPM_PARTITION_CONFIG_INIT_C,
    partitionStat  => XPM_PARTITION_STATUS_INIT_C,
    pllCfg         => XPM_PLL_CONFIG_INIT_C,
    pllStat        => XPM_PLL_STATUS_INIT_C,
    inhibitCfg     => XPM_INHIBIT_CONFIG_INIT_C,
    axilReadSlave  => AXI_LITE_READ_SLAVE_INIT_C,
    axilWriteSlave => AXI_LITE_WRITE_SLAVE_INIT_C,
    axilRdEn       => (others=>'1'),
    linkDebug      => (others=>'0'),
    tagStream      => '0',
    anaWrCount     => (others=>(others=>'0')));

  constant TAG_AXIS_CONFIG_C : AxiStreamConfigType := ssiAxiStreamConfig(8);
  signal tagMaster : AxiStreamMasterType;
  
  signal r    : RegType := REG_INIT_C;
  signal r_in : RegType;

  signal pll_stat    : slv(2*NAmcs-1 downto 0);
  signal pllStat     : slv(2*NAmcs-1 downto 0);
  signal pllCount    : SlVectorArray(2*NAmcs-1 downto 0, 2 downto 0);

  type AnaRdArray is array (natural range<>) of SlVectorArray(0 downto 0,31 downto 0);
  signal anaRdCount  : AnaRdArray(NPartitions-1 downto 0);
  
  signal s    : XpmStatusType;
  signal sbpLinkUp : slv(NBPLinks downto 0);
  
begin

  dbgChan        <= r.linkDebug(dbgChan'range);
  config         <= r.config;
  axilReadSlave  <= r.axilReadSlave;
  axilWriteSlave <= r.axilWriteSlave;
  axilUpdate     <= r.axilRdEn;

  --
  --  Still need to cross clock-domains for register readout of:
  --    link status (32 links)
  --    partition inhibit counts (from 32 links for each partition)
  --
  
  GEN_BPLINK : entity work.SynchronizerVector
    generic map ( WIDTH_G => sbpLinkUp'length )
    port map ( clk     => regClk,
               dataIn  => status.bpLinkUp,
               dataOut => sbpLinkUp );
  
  GEN_PART : for i in 0 to NPartitions-1 generate
    U_Sync64_ena : entity work.SynchronizerFifo
      generic map ( DATA_WIDTH_G => 64 )
      port map ( wr_clk => staClk, rd_clk=> axilClk, rd_en=> r.axilRdEn(i),
                 din  => status.partition(i).l0Select.enabled  ,
                 dout => s.partition(i).l0Select.enabled);
    U_Sync64_inh : entity work.SynchronizerFifo
      generic map ( DATA_WIDTH_G => 64 )
      port map ( wr_clk => staClk, rd_clk=> axilClk, rd_en=> r.axilRdEn(i),
                 din  => status.partition(i).l0Select.inhibited  ,
                 dout => s.partition(i).l0Select.inhibited);
    U_Sync64_num : entity work.SynchronizerFifo
      generic map ( DATA_WIDTH_G => 64 )
      port map ( wr_clk => staClk, rd_clk=> axilClk, rd_en=> r.axilRdEn(i),
                 din  => status.partition(i).l0Select.num  ,
                 dout => s.partition(i).l0Select.num);
    U_Sync64_nin : entity work.SynchronizerFifo
      generic map ( DATA_WIDTH_G => 64 )
      port map ( wr_clk => staClk, rd_clk=> axilClk, rd_en=> r.axilRdEn(i),
                 din  => status.partition(i).l0Select.numInh  ,
                 dout => s.partition(i).l0Select.numInh);
    U_Sync64_nac : entity work.SynchronizerFifo
      generic map ( DATA_WIDTH_G => 64 )
      port map ( wr_clk => staClk, rd_clk=> axilClk, rd_en=> r.axilRdEn(i),
                 din  => status.partition(i).l0Select.numAcc  ,
                 dout => s.partition(i).l0Select.numAcc);
    U_SyncAna : entity work.SyncStatusVector
      generic map ( WIDTH_G     => 1,
                    CNT_WIDTH_G => 32 )
      port map ( statusIn  => status.partition(i).anaRd(1 downto 1),
                 statusOut => open,
                 cntRstIn  => r.config.partition(i).analysis.rst(1),
                 rollOverEnIn => (others=>'1'),
                 cntOut    => anaRdCount(i),
                 wrClk     => staClk,
                 rdClk     => axilClk );
  end generate;
  
  GEN_LOL : for i in 0 to NAmcs-1 generate
    pll_stat(2*i+0) <= pllStatus(i).los;
    pll_stat(2*i+1) <= pllStatus(i).lol;
  end generate;
    
  U_StatLol : entity work.SyncStatusVector
     generic map ( COMMON_CLK_G => true,
                   WIDTH_G      => 2*NAmcs,
                   CNT_WIDTH_G  => 3 )
     port map ( statusIn  => pll_stat,
                statusOut => pllStat,
                cntRstIn  => '0',
                rollOverEnIn => (others=>'1'),
                cntOut    => pllCount,
                wrClk     => axilClk,
                rdClk     => axilClk );
                
  U_AnalysisFifo : entity work.AxiStreamFifo
    generic map ( SLAVE_AXI_CONFIG_G  => ETH_AXIS_CONFIG_C,
                  MASTER_AXI_CONFIG_G => TAG_AXIS_CONFIG_C )
    port map ( sAxisClk     => axilClk,
               sAxisRst     => axilRst,
               sAxisMaster  => ibDebugMaster,
               sAxisSlave   => ibDebugSlave,
               mAxisClk     => axilClk,
               mAxisRst     => axilRst,
               mAxisMaster  => tagMaster,
               mAxisSlave   => r_in.tagSlave );

  comb : process (r, axilReadMaster, axilWriteMaster, tagMaster, status, s, axilRst,
                  pllStatus, pllCount, pllStat, anaRdCount, sbpLinkUp) is
    variable v          : RegType;
    variable axilStatus : AxiLiteStatusType;
    variable ip         : integer;
    variable il         : integer;
    variable ia         : integer;
    -- Shorthand procedures for read/write register
    procedure axilRegRW(addr : in slv; offset : in integer; reg : inout slv) is
    begin
      axiSlaveRegister(axilWriteMaster, axilReadMaster,
                       v.axilWriteSlave, v.axilReadSlave, axilStatus,
                       addr, offset, reg, false, "0");
    end procedure;
    procedure axilRegRW(addr : in slv; offset : in integer; reg : inout sl) is
    begin
      axiSlaveRegister(axilWriteMaster, axilReadMaster,
                       v.axilWriteSlave, v.axilReadSlave, axilStatus,
                       addr, offset, reg, false, '0');
    end procedure;
    -- Shorthand procedures for read only registers
    procedure axilRegR (addr : in slv; offset : in integer; reg : in slv) is
    begin
      axiSlaveRegister(axilReadMaster, v.axilReadSlave, axilStatus,
                       addr, offset, reg);
    end procedure;
    procedure axilRegR (addr : in slv; offset : in integer; reg : in sl) is
    begin
      axiSlaveRegister(axilReadMaster, v.axilReadSlave, axilStatus,
                       addr, offset, reg);
    end procedure;
    procedure axilRegR64 (addr : in slv; reg : in slv) is
    begin
      axilRegR(addr+0,0,reg(31 downto  0));
      axilRegR(addr+4,0,reg(63 downto 32));
    end procedure;
  begin
    v := r;
    -- reset strobing signals
    v.axilReadSlave.rdata := (others=>'0');
    v.partitionCfg.message.insert := '0';
    v.tagSlave.tReady      := '1';

    ip := conv_integer(r.partition);
    il := conv_integer(r.link(3 downto 0));
    ia := conv_integer(r.amc);
    
    if r.load='1' then
      if r.link(4)='0' then
        v.linkCfg      := r.config.dsLink(il);
      else
        v.linkCfg      := r.config.bpLink(il);
      end if;
      v.partitionCfg := r.config.partition(ip);
      v.pllCfg       := r.config.pll      (ia);
    else
      if r.link(4)='0' then
        v.config.dsLink (il)      := r.linkCfg;
      else
        v.config.bpLink (il)      := r.linkCfg;
      end if;
      v.config.partition(ip)      := r.partitionCfg;
      v.config.pll      (ia)      := r.pllCfg;
    end if;

    if r.link(4)='0' then
      v.linkStat         := status.dsLink (il);
    elsif r.link(3 downto 0)=toSlv(NBPLinks,4) then
      v.linkStat         := XPM_LINK_STATUS_INIT_C;
      v.linkStat.txReady := sbpLinkUp(il);
    else
      v.linkStat         := XPM_LINK_STATUS_INIT_C;
      v.linkStat.rxReady := sbpLinkUp(il);
    end if;
    v.partitionStat := status.partition(ip);
    v.pllStat       := pllStatus       (ia);
    
    -- Determine the transaction type
    axiSlaveWaitTxn(axilWriteMaster, axilReadMaster, v.axilWriteSlave, v.axilReadSlave, axilStatus);
    v.axilReadSlave.rdata := (others=>'0');
    
    -- Read/write to the configuration registers
    -- Read only from status registers

    axilRegR  (toSlv(  0,12),  0, status.paddr);
    axilRegRW (toSlv(  4,12),  0, v.partition);
    axilRegRW (toSlv(  4,12),  4, v.link);
    axilRegRW (toSlv(  4,12), 10, v.linkDebug);
    axilRegRW (toSlv(  4,12), 16, v.amc);
    axilRegRW (toSlv(  4,12), 20, v.inhibit);
    axilRegRW (toSlv(  4,12), 24, v.tagStream);
    
    v.load := '0';
    v.linkCfg.txDelayRst   := '0';

    if axilStatus.writeEnable='1' then
      if std_match(axilWriteMaster.awaddr(11 downto 0),toSlv(4,12)) then
        v.load := '1';
      end if;
        
      if std_match(axilWriteMaster.awaddr(11 downto 0),toSlv(8,12)) then
        v.linkCfg.txDelayRst := '1';
      end if;
    end if;
    
    axilRegRW(toSlv(8,12),    0, v.linkCfg.txDelay);
    axilRegRW(toSlv(8,12),   20, v.linkCfg.partition);
    axilRegRW(toSlv(8,12),   24, v.linkCfg.trigsrc);
    axilRegRW(toSlv(8,12),   28, v.linkCfg.loopback);
    axilRegRW(toSlv(8,12),   29, v.linkCfg.txReset);
    axilRegRW(toSlv(8,12),   30, v.linkCfg.rxReset);
    axilRegRW(toSlv(8,12),   31, v.linkCfg.enable);
    
    axilRegR (toSlv(12,12),   0, r.linkStat.rxErrCnts);
    axilRegR (toSlv(12,12),  16, r.linkStat.txResetDone);
    axilRegR (toSlv(12,12),  17, r.linkStat.txReady);
    axilRegR (toSlv(12,12),  18, r.linkStat.rxResetDone);
    axilRegR (toSlv(12,12),  19, r.linkStat.rxReady);
    axilRegR (toSlv(12,12),  20, r.linkStat.rxIsXpm);

    axilRegRW(toSlv(16,12),  0, v.pllCfg.bwSel);
    axilRegRW(toSlv(16,12),  4, v.pllCfg.frqTbl);
    axilRegRW(toSlv(16,12),  8, v.pllCfg.frqSel);
    axilRegRW(toSlv(16,12), 16, v.pllCfg.rate);
    axilRegRW(toSlv(16,12), 20, v.pllCfg.inc);
    axilRegRW(toSlv(16,12), 21, v.pllCfg.dec);
    axilRegRW(toSlv(16,12), 22, v.pllCfg.bypass);
    axilRegRW(toSlv(16,12), 23, v.pllCfg.rstn);
    axilRegR (toSlv(16,12), 24, muxSlVectorArray( pllCount, 2*ia+0));
    axilRegR (toSlv(16,12), 27, pllStat(2*ia+0));
    axilRegR (toSlv(16,12), 28, muxSlVectorArray( pllCount, 2*ia+1));
    axilRegR (toSlv(16,12), 31, pllStat(2*ia+1));

    axilRegRW (toSlv(20,12), 0, v.partitionCfg.l0Select.reset);
    axilRegRW (toSlv(20,12),16, v.partitionCfg.l0Select.enabled);
    axilRegRW (toSlv(20,12),31, v.axilRdEn(ip));
    axilRegRW (toSlv(24,12), 0, v.partitionCfg.l0Select.rateSel);
    axilRegRW (toSlv(24,12),16, v.partitionCfg.l0Select.destSel);

    axilRegR64(toSlv(28,12), s.partition(ip).l0Select.enabled);
    axilRegR64(toSlv(36,12), s.partition(ip).l0Select.inhibited);
    axilRegR64(toSlv(44,12), s.partition(ip).l0Select.num);
    axilRegR64(toSlv(52,12), s.partition(ip).l0Select.numInh);
    axilRegR64(toSlv(60,12), s.partition(ip).l0Select.numAcc);
    axilRegR64(toSlv(68,12), s.partition(ip).l1Select.numAcc);

    axilRegRW (toSlv(76,12),  0, v.partitionCfg.l1Select.clear);
    axilRegRW (toSlv(76,12), 16, v.partitionCfg.l1Select.enable);
    axilRegRW (toSlv(80,12),  0, v.partitionCfg.l1Select.trigsrc);
    axilRegRW (toSlv(80,12),  4, v.partitionCfg.l1Select.trigword);
    axilRegRW (toSlv(80,12), 16, v.partitionCfg.l1Select.trigwr);
      
    axilRegRW (toSlv(84,12), 0, v.partitionCfg.analysis.rst);
    axilRegRW (toSlv(88,12), 0, v.partitionCfg.analysis.tag);
    axilRegRW (toSlv(92,12), 0, v.partitionCfg.analysis.push);
    axilRegR  (toSlv(96,12), 0, r.anaWrCount(ip));
    axilRegR  (toSlv(100,12), 0, muxSlVectorArray( anaRdCount(ip), 0));

    axilRegRW (toSlv(104,12), 0, v.partitionCfg.pipeline.depth);

    axilRegRW (toSlv(108,12),15, v.partitionCfg.message.insert);
    axilRegRW (toSlv(108,12), 0, v.partitionCfg.message.hdr);
    axilRegRW (toSlv(112,12), 0, v.partitionCfg.message.payload);

    for j in r.partitionCfg.inhibit.setup'range loop
      axilRegRW (toSlv(128+j*4,12),  0, v.partitionCfg.inhibit.setup(j).interval);
      axilRegRW (toSlv(128+j*4,12), 12, v.partitionCfg.inhibit.setup(j).limit);
      axilRegRW (toSlv(128+j*4,12), 31, v.partitionCfg.inhibit.setup(j).enable);
    end loop;

    for j in 0 to 31 loop
      axilRegR (toSlv(144+j*4,12), 0, r.partitionStat.inhibit.counts(j));
    end loop;

    if r.partitionCfg.analysis.rst(1)='1' then
      v.anaWrCount(ip) := (others=>'0');
    elsif r.partitionCfg.analysis.push(1)='1' then
      v.anaWrCount(ip) := r.anaWrCount(ip)+1;
    end if;
      
    if r.config.tagstream='0' then
      v.tagSlave.tReady := '0';
    elsif tagMaster.tValid='1' then
      ip := conv_integer(tagMaster.tDest(3 downto 0));
      v.config.partition(ip).analysis.tag  := tagMaster.tData(31 downto  0);
      v.config.partition(ip).analysis.push := tagMaster.tData(35 downto 34);
    end if;

    -- Set the status
    axiSlaveDefault(axilWriteMaster, axilReadMaster, v.axilWriteSlave, v.axilReadSlave, axilStatus, AXI_RESP_OK_C);

    ----------------------------------------------------------------------------------------------
    -- Reset
    ----------------------------------------------------------------------------------------------
    if (axilRst = '1') then
      v := REG_INIT_C;
    end if;

    r_in <= v;
  end process;

  seq : process (axilClk) is
  begin
    if rising_edge(axilClk) then
      r <= r_in;
    end if;
  end process;
end rtl;
